//Verilog HDL for "BioZ_EMG_Model", "BioZ_SIGGEN_DACCtrl" "functional"


module BioZ_SigGen_DACCtrl_2 (
CountEnable,
Clk,
Clk_IF,
Resetn,
StepNum,
P,
clk_IF_P,
clk_IF_N,
clk_merged_IP,
clk_merged_IN,
clk_merged_QP,
clk_merged_QN,
IP,
IN,
QP,
QN
);


//Inputs
input CountEnable;
input Clk;
input Clk_IF;
input Resetn;
input StepNum;


//Outputs
//output wire P1,P2,P3,P4,P5; //Control signals for the DAC
output reg [32:0] P; //Control signals for the DAC
output wire IP,IN; // in-phase (I) reference clock
output wire QP,QN; // quadrature (Q) reference clock
output wire clk_IF_P, clk_IF_N; // IF reference clock
output wire clk_merged_IP,clk_merged_IN, clk_merged_QP,clk_merged_QN; // I/Q merged clocks (I/Q XNOR IF)

reg [32:0] S64;
reg [32:0] S32;
reg [32:0] S16;

reg [5:0] count;
reg [5:0] count_IF;

reg IP_aux, QP_aux, IN_aux, QN_aux, IF_P_aux, IF_N_aux, Q_samp;

// 5bit counter state machine
always @(posedge Clk, negedge Resetn)
begin
    if (Resetn == 0) begin
        count <= 0;
    end else begin
        count <= count + 1;    
    end    
end

always @(posedge Clk_IF, negedge Resetn)
begin
    if (Resetn == 0) begin
        count_IF <= 0;
    end else begin
        count_IF <= count_IF + 1;    
    end    
end

// AMS VERSION 32 steps - 16 steps

//Intermediate signals 64 steps
always @(CountEnable, count)
begin
    if (CountEnable == 1) begin
        case(count)
            0:  S64 = 33'b0_0000_0000_0000_0000_0000_0000_0000_0001; //0 0V         
            1:  S64 = 33'b0_0000_0000_0000_0000_0000_0000_0000_0010;
            2:  S64 = 33'b0_0000_0000_0000_0000_0000_0000_0000_0100;
            3:  S64 = 33'b0_0000_0000_0000_0000_0000_0000_0000_1000;
            4:  S64 = 33'b0_0000_0000_0000_0000_0000_0000_0001_0000;
            5:  S64 = 33'b0_0000_0000_0000_0000_0000_0000_0010_0000;
            6:  S64 = 33'b0_0000_0000_0000_0000_0000_0000_0100_0000;
            7:  S64 = 33'b0_0000_0000_0000_0000_0000_0000_1000_0000;
            8:  S64 = 33'b0_0000_0000_0000_0000_0000_0001_0000_0000; //8 +0.5V
            9:  S64 = 33'b0_0000_0000_0000_0000_0000_0010_0000_0000;
            10: S64 = 33'b0_0000_0000_0000_0000_0000_0100_0000_0000;
            11: S64 = 33'b0_0000_0000_0000_0000_0000_1000_0000_0000;
            12: S64 = 33'b0_0000_0000_0000_0000_0001_0000_0000_0000;
            13: S64 = 33'b0_0000_0000_0000_0000_0010_0000_0000_0000;
            14: S64 = 33'b0_0000_0000_0000_0000_0100_0000_0000_0000;
            15: S64 = 33'b0_0000_0000_0000_0000_1000_0000_0000_0000;
            16: S64 = 33'b0_0000_0000_0000_0001_0000_0000_0000_0000; //16 +1V
            17: S64 = 33'b0_0000_0000_0000_0000_1000_0000_0000_0000;
            18: S64 = 33'b0_0000_0000_0000_0000_0100_0000_0000_0000;
            19: S64 = 33'b0_0000_0000_0000_0000_0010_0000_0000_0000;
            20: S64 = 33'b0_0000_0000_0000_0000_0001_0000_0000_0000;
            21: S64 = 33'b0_0000_0000_0000_0000_0000_1000_0000_0000;
            22: S64 = 33'b0_0000_0000_0000_0000_0000_0100_0000_0000;
            23: S64 = 33'b0_0000_0000_0000_0000_0000_0010_0000_0000;
            24: S64 = 33'b0_0000_0000_0000_0000_0000_0001_0000_0000; //8 +0.5V
            25: S64 = 33'b0_0000_0000_0000_0000_0000_0000_1000_0000;
            26: S64 = 33'b0_0000_0000_0000_0000_0000_0000_0100_0000;
            27: S64 = 33'b0_0000_0000_0000_0000_0000_0000_0010_0000;
            28: S64 = 33'b0_0000_0000_0000_0000_0000_0000_0001_0000;
            29: S64 = 33'b0_0000_0000_0000_0000_0000_0000_0000_1000;
            30: S64 = 33'b0_0000_0000_0000_0000_0000_0000_0000_0100;
            31: S64 = 33'b0_0000_0000_0000_0000_0000_0000_0000_0010;
            32: S64 = 33'b0_0000_0000_0000_0000_0000_0000_0000_0001; //0 0V     
            33: S64 = 33'b0_0000_0000_0000_0010_0000_0000_0000_0000;
            34: S64 = 33'b0_0000_0000_0000_0100_0000_0000_0000_0000;
            35: S64 = 33'b0_0000_0000_0000_1000_0000_0000_0000_0000;
            36: S64 = 33'b0_0000_0000_0001_0000_0000_0000_0000_0000;
            37: S64 = 33'b0_0000_0000_0010_0000_0000_0000_0000_0000;
            38: S64 = 33'b0_0000_0000_0100_0000_0000_0000_0000_0000;
            39: S64 = 33'b0_0000_0000_1000_0000_0000_0000_0000_0000;
            40: S64 = 33'b0_0000_0001_0000_0000_0000_0000_0000_0000; //32 -0.5V
            41: S64 = 33'b0_0000_0010_0000_0000_0000_0000_0000_0000;
            42: S64 = 33'b0_0000_0100_0000_0000_0000_0000_0000_0000;
            43: S64 = 33'b0_0000_1000_0000_0000_0000_0000_0000_0000;
            44: S64 = 33'b0_0001_0000_0000_0000_0000_0000_0000_0000;
            45: S64 = 33'b0_0010_0000_0000_0000_0000_0000_0000_0000;
            46: S64 = 33'b0_0100_0000_0000_0000_0000_0000_0000_0000;
            47: S64 = 33'b0_1000_0000_0000_0000_0000_0000_0000_0000;
            48: S64 = 33'b1_0000_0000_0000_0000_0000_0000_0000_0000; //64 -1V
            49: S64 = 33'b0_1000_0000_0000_0000_0000_0000_0000_0000;
            50: S64 = 33'b0_0100_0000_0000_0000_0000_0000_0000_0000;
            51: S64 = 33'b0_0010_0000_0000_0000_0000_0000_0000_0000;
            52: S64 = 33'b0_0001_0000_0000_0000_0000_0000_0000_0000;
            53: S64 = 33'b0_0000_1000_0000_0000_0000_0000_0000_0000;
            54: S64 = 33'b0_0000_0100_0000_0000_0000_0000_0000_0000;
            55: S64 = 33'b0_0000_0010_0000_0000_0000_0000_0000_0000;
            56: S64 = 33'b0_0000_0001_0000_0000_0000_0000_0000_0000; //32 -0.5V
            57: S64 = 33'b0_0000_0000_1000_0000_0000_0000_0000_0000;
            58: S64 = 33'b0_0000_0000_0100_0000_0000_0000_0000_0000;
            59: S64 = 33'b0_0000_0000_0010_0000_0000_0000_0000_0000;
            60: S64 = 33'b0_0000_0000_0001_0000_0000_0000_0000_0000;
            61: S64 = 33'b0_0000_0000_0000_1000_0000_0000_0000_0000;
            62: S64 = 33'b0_0000_0000_0000_0100_0000_0000_0000_0000;
            63: S64 = 33'b0_0000_0000_0000_0010_0000_0000_0000_0000;
            default: S64 = 33'b0_0000_0000_0000_0000_0000_0000_0000_0001; //0 0V    
         endcase   
    end else begin
            S64 = 33'b0_0000_0000_0000_0000_0000_0000_0000_0001; //0 0V  
    end
end


//Intermediate signals 32 steps
always @(CountEnable, count)
begin
    if (CountEnable == 1) begin
        case(count)
            0:  S32 = 33'b0_0000_0000_0000_0000_0000_0000_0000_0001; //0 0V         
            1:  S32 = 33'b0_0000_0000_0000_0000_0000_0000_0000_0100;
            2:  S32 = 33'b0_0000_0000_0000_0000_0000_0000_0001_0000;
            3:  S32 = 33'b0_0000_0000_0000_0000_0000_0000_0100_0000;
            4:  S32 = 33'b0_0000_0000_0000_0000_0000_0001_0000_0000; //8 +0.5V
            5:  S32 = 33'b0_0000_0000_0000_0000_0000_0100_0000_0000;
            6:  S32 = 33'b0_0000_0000_0000_0000_0001_0000_0000_0000;
            7:  S32 = 33'b0_0000_0000_0000_0000_0100_0000_0000_0000;
            8:  S32 = 33'b0_0000_0000_0000_0001_0000_0000_0000_0000; //16 +1V
            9:  S32 = 33'b0_0000_0000_0000_0000_0100_0000_0000_0000;
            10: S32 = 33'b0_0000_0000_0000_0000_0001_0000_0000_0000;
            11: S32 = 33'b0_0000_0000_0000_0000_0000_0100_0000_0000;
            12: S32 = 33'b0_0000_0000_0000_0000_0000_0001_0000_0000; //8 +0.5V
            13: S32 = 33'b0_0000_0000_0000_0000_0000_0000_0100_0000;
            14: S32 = 33'b0_0000_0000_0000_0000_0000_0000_0001_0000;
            15: S32 = 33'b0_0000_0000_0000_0000_0000_0000_0000_0100;
            16: S32 = 33'b0_0000_0000_0000_0000_0000_0000_0000_0001; //0 0V
            17: S32 = 33'b0_0000_0000_0000_0100_0000_0000_0000_0000;
            18: S32 = 33'b0_0000_0000_0001_0000_0000_0000_0000_0000;
            19: S32 = 33'b0_0000_0000_0100_0000_0000_0000_0000_0000;
            20: S32 = 33'b0_0000_0001_0000_0000_0000_0000_0000_0000; //32 -0.5V
            21: S32 = 33'b0_0000_0100_0000_0000_0000_0000_0000_0000;
            22: S32 = 33'b0_0001_0000_0000_0000_0000_0000_0000_0000;
            23: S32 = 33'b0_0100_0000_0000_0000_0000_0000_0000_0000;
            24: S32 = 33'b1_0000_0000_0000_0000_0000_0000_0000_0000; //64 -1V
            25: S32 = 33'b0_0100_0000_0000_0000_0000_0000_0000_0000;
            26: S32 = 33'b0_0001_0000_0000_0000_0000_0000_0000_0000;
            27: S32 = 33'b0_0000_0100_0000_0000_0000_0000_0000_0000;
            28: S32 = 33'b0_0000_0001_0000_0000_0000_0000_0000_0000; //32 -0.5V
            29: S32 = 33'b0_0000_0000_0100_0000_0000_0000_0000_0000;
            30: S32 = 33'b0_0000_0000_0001_0000_0000_0000_0000_0000;
            31: S32 = 33'b0_0000_0000_0000_0100_0000_0000_0000_0000;
            32: S32 = 33'b0_0000_0000_0000_0000_0000_0000_0000_0001; //0 0V     
            33: S32 = 33'b0_0000_0000_0000_0000_0000_0000_0000_0100;
            34: S32 = 33'b0_0000_0000_0000_0000_0000_0000_0001_0000;
            35: S32 = 33'b0_0000_0000_0000_0000_0000_0000_0100_0000;
            36: S32 = 33'b0_0000_0000_0000_0000_0000_0001_0000_0000; //8 +0.5V
            37: S32 = 33'b0_0000_0000_0000_0000_0000_0100_0000_0000;
            38: S32 = 33'b0_0000_0000_0000_0000_0001_0000_0000_0000;
            39: S32 = 33'b0_0000_0000_0000_0000_0100_0000_0000_0000;
            40: S32 = 33'b0_0000_0000_0000_0001_0000_0000_0000_0000; //16 +1V
            41: S32 = 33'b0_0000_0000_0000_0000_0100_0000_0000_0000;
            42: S32 = 33'b0_0000_0000_0000_0000_0001_0000_0000_0000;
            43: S32 = 33'b0_0000_0000_0000_0000_0000_0100_0000_0000;
            44: S32 = 33'b0_0000_0000_0000_0000_0000_0001_0000_0000; //8 +0.5V
            45: S32 = 33'b0_0000_0000_0000_0000_0000_0000_0100_0000;
            46: S32 = 33'b0_0000_0000_0000_0000_0000_0000_0001_0000;
            47: S32 = 33'b0_0000_0000_0000_0000_0000_0000_0000_0100;
            48: S32 = 33'b0_0000_0000_0000_0000_0000_0000_0000_0001; //0 0V  
            49: S32 = 33'b0_0000_0000_0000_0100_0000_0000_0000_0000;
            50: S32 = 33'b0_0000_0000_0001_0000_0000_0000_0000_0000;
            51: S32 = 33'b0_0000_0000_0100_0000_0000_0000_0000_0000;
            52: S32 = 33'b0_0000_0001_0000_0000_0000_0000_0000_0000; //32 -0.5V
            53: S32 = 33'b0_0000_0100_0000_0000_0000_0000_0000_0000;
            54: S32 = 33'b0_0001_0000_0000_0000_0000_0000_0000_0000;
            55: S32 = 33'b0_0100_0000_0000_0000_0000_0000_0000_0000;
            56: S32 = 33'b1_0000_0000_0000_0000_0000_0000_0000_0000; //64 -1V
            57: S32 = 33'b0_0100_0000_0000_0000_0000_0000_0000_0000;
            58: S32 = 33'b0_0001_0000_0000_0000_0000_0000_0000_0000;
            59: S32 = 33'b0_0000_0100_0000_0000_0000_0000_0000_0000;
            60: S32 = 33'b0_0000_0001_0000_0000_0000_0000_0000_0000; //32 -0.5V
            61: S32 = 33'b0_0000_0000_0100_0000_0000_0000_0000_0000;
            62: S32 = 33'b0_0000_0000_0001_0000_0000_0000_0000_0000;
            63: S32 = 33'b0_0000_0000_0000_0100_0000_0000_0000_0000;
            default: S32 = 33'b0_0000_0000_0000_0000_0000_0000_0000_0001; //0 0V 
         endcase   
    end else begin
            S32 = 33'b0_0000_0000_0000_0000_0000_0000_0000_0001; //0 0V  
    end
end

//Intermediate signals 16 steps
always @(CountEnable, count)
begin
    if (CountEnable == 1) begin
        case(count)
            0:  S16 = 33'b0_0000_0000_0000_0000_0000_0000_0000_0001; //0 0V         
            1:  S16 = 33'b0_0000_0000_0000_0000_0000_0000_0001_0000;
            2:  S16 = 33'b0_0000_0000_0000_0000_0000_0001_0000_0000;
            3:  S16 = 33'b0_0000_0000_0000_0000_0001_0000_0000_0000;
            4:  S16 = 33'b0_0000_0000_0000_0001_0000_0000_0000_0000; //8 +0.5V
            5:  S16 = 33'b0_0000_0000_0000_0000_0001_0000_0000_0000;
            6:  S16 = 33'b0_0000_0000_0000_0000_0000_0001_0000_0000;
            7:  S16 = 33'b0_0000_0000_0000_0000_0000_0000_0001_0000;
            8:  S16 = 33'b0_0000_0000_0000_0000_0000_0000_0000_0001; //16 +1V
            9:  S16 = 33'b0_0000_0000_0001_0000_0000_0000_0000_0000;
            10: S16 = 33'b0_0000_0001_0000_0000_0000_0000_0000_0000;
            11: S16 = 33'b0_0001_0000_0000_0000_0000_0000_0000_0000;
            12: S16 = 33'b1_0000_0000_0000_0000_0000_0000_0000_0000; //8 +0.5V
            13: S16 = 33'b0_0001_0000_0000_0000_0000_0000_0000_0000;
            14: S16 = 33'b0_0000_0001_0000_0000_0000_0000_0000_0000;
            15: S16 = 33'b0_0000_0000_0001_0000_0000_0000_0000_0000;
            16: S16 = 33'b0_0000_0000_0000_0000_0000_0000_0000_0001; //0 0V
            17: S16 = 33'b0_0000_0000_0000_0000_0000_0000_0001_0000;
            18: S16 = 33'b0_0000_0000_0000_0000_0000_0001_0000_0000;
            19: S16 = 33'b0_0000_0000_0000_0000_0001_0000_0000_0000;
            20: S16 = 33'b0_0000_0000_0000_0001_0000_0000_0000_0000; //32 -0.5V
            21: S16 = 33'b0_0000_0000_0000_0000_0001_0000_0000_0000;
            22: S16 = 33'b0_0000_0000_0000_0000_0000_0001_0000_0000;
            23: S16 = 33'b0_0000_0000_0000_0000_0000_0000_0001_0000;
            24: S16 = 33'b0_0000_0000_0000_0000_0000_0000_0000_0001; //64 -1V
            25: S16 = 33'b0_0000_0000_0001_0000_0000_0000_0000_0000;
            26: S16 = 33'b0_0000_0001_0000_0000_0000_0000_0000_0000;
            27: S16 = 33'b0_0001_0000_0000_0000_0000_0000_0000_0000;
            28: S16 = 33'b1_0000_0000_0000_0000_0000_0000_0000_0000; //32 -0.5V
            29: S16 = 33'b0_0001_0000_0000_0000_0000_0000_0000_0000;
            30: S16 = 33'b0_0000_0001_0000_0000_0000_0000_0000_0000;
            31: S16 = 33'b0_0000_0000_0001_0000_0000_0000_0000_0000;
            32: S16 = 33'b0_0000_0000_0000_0000_0000_0000_0000_0001; //0 0V     
            33: S16 = 33'b0_0000_0000_0000_0000_0000_0000_0001_0000;
            34: S16 = 33'b0_0000_0000_0000_0000_0000_0001_0000_0000;
            35: S16 = 33'b0_0000_0000_0000_0000_0001_0000_0000_0000;
            36: S16 = 33'b0_0000_0000_0000_0001_0000_0000_0000_0000; //8 +0.5V
            37: S16 = 33'b0_0000_0000_0000_0000_0001_0000_0000_0000;
            38: S16 = 33'b0_0000_0000_0000_0000_0000_0001_0000_0000;
            39: S16 = 33'b0_0000_0000_0000_0000_0000_0000_0001_0000;
            40: S16 = 33'b0_0000_0000_0000_0000_0000_0000_0000_0001; //16 +1V
            41: S16 = 33'b0_0000_0000_0001_0000_0000_0000_0000_0000;
            42: S16 = 33'b0_0000_0001_0000_0000_0000_0000_0000_0000;
            43: S16 = 33'b0_0001_0000_0000_0000_0000_0000_0000_0000;
            44: S16 = 33'b1_0000_0000_0000_0000_0000_0000_0000_0000; //8 +0.5V
            45: S16 = 33'b0_0001_0000_0000_0000_0000_0000_0000_0000;
            46: S16 = 33'b0_0000_0001_0000_0000_0000_0000_0000_0000;
            47: S16 = 33'b0_0000_0000_0001_0000_0000_0000_0000_0000;
            48: S16 = 33'b0_0000_0000_0000_0000_0000_0000_0000_0001; //0 0V  
            49: S16 = 33'b0_0000_0000_0000_0000_0000_0000_0001_0000;
            50: S16 = 33'b0_0000_0000_0000_0000_0000_0001_0000_0000;
            51: S16 = 33'b0_0000_0000_0000_0000_0001_0000_0000_0000;
            52: S16 = 33'b0_0000_0000_0000_0001_0000_0000_0000_0000; //32 -0.5V
            53: S16 = 33'b0_0000_0000_0000_0000_0001_0000_0000_0000;
            54: S16 = 33'b0_0000_0000_0000_0000_0000_0001_0000_0000;
            55: S16 = 33'b0_0000_0000_0000_0000_0000_0000_0001_0000;
            56: S16 = 33'b0_0000_0000_0000_0000_0000_0000_0000_0001; //64 -1V
            57: S16 = 33'b0_0000_0000_0001_0000_0000_0000_0000_0000;
            58: S16 = 33'b0_0000_0001_0000_0000_0000_0000_0000_0000;
            59: S16 = 33'b0_0001_0000_0000_0000_0000_0000_0000_0000;
            60: S16 = 33'b1_0000_0000_0000_0000_0000_0000_0000_0000; //32 -0.5V
            61: S16 = 33'b0_0001_0000_0000_0000_0000_0000_0000_0000;
            62: S16 = 33'b0_0000_0001_0000_0000_0000_0000_0000_0000;
            63: S16 = 33'b0_0000_0000_0001_0000_0000_0000_0000_0000;
            default: S16 = 33'b0_0000_0000_0000_0000_0000_0000_0000_0001; //0 0V 
         endcase   
    end else begin
            S16 = 33'b0_0000_0000_0000_0000_0000_0000_0000_0001; //0 0V  
    end
end

always @(StepNum,S16,S32,S64)
begin
	case(StepNum) // 00 selects 64 steps, 01 selects 32 steps, 10 selects 16 steps
		2'b00: P = S64;
		2'b01: P = S32;
		2'b10: P = S16;
		default:  P = S64;
    endcase
end

// IF Outputs


always @(StepNum,count_IF)
begin
	case(StepNum) // 00 selects 64 steps, 01 selects 32 steps, 10 selects 16 steps
		2'b00: begin
			IF_P_aux <= ~count_IF[5];
			IF_N_aux <= count_IF[5];
		end
		2'b01: begin // 32 Steps
			IF_P_aux <= ~count_IF[4];
			IF_N_aux <= count_IF[4];
		end
		2'b10: begin // 16 steps
			IF_P_aux <= ~count_IF[3];
			IF_N_aux <= count_IF[3];
		end
		default: begin
			IF_P_aux <= ~count_IF[5];
			IF_N_aux <= count_IF[5];
		end
    endcase
end

assign clk_IF_P = IF_P_aux;
assign clk_IF_N = IF_N_aux;

// I/Q Outputs

always @(StepNum,count)
begin
	if(StepNum == 0) begin // 32 Steps
		IP_aux <= ~count[4];
		IN_aux <= count[4];	
	end else begin // 16 steps
		IP_aux <= ~count[3];
		IN_aux <= count[3];	
	end
end

assign IP = IP_aux;
assign IN = IN_aux;

//always @(StepNum,count)
//begin
//	if(StepNum == 0) begin //32 steps
//		QP_aux = ~count[4];
//		QN_aux <= count[4];	
//	end else begin //16 steps
//		QP_aux = ~count[3];
//		QN_aux <= count[3];	
//	end
//end

//assign QP = QP_aux;
//assign QN = QN_aux;

// clk_merged Outputs

assign clk_merged_IP = (IP ~^ clk_IF_P);
assign clk_merged_IN = ~clk_merged_IP;
assign clk_merged_QP = (QP ~^ clk_IF_P);
assign clk_merged_QN = ~clk_merged_QP;

//Q is created by sampling I exactly in the middle of the high pulse. 
//Aux_Q is the clock used to sample I;

always @(StepNum,count)
begin
    if(StepNum == 0) begin //32 steps
        Q_samp = count[3];
    end else begin //16 steps
        Q_samp = count[2];
    end
end

always @(posedge Q_samp, negedge Resetn)
begin
	if (Resetn == 0) begin
		QP_aux <= 0;
	end else begin
		QP_aux <= IP;
	end    
end

assign QP = QP_aux;
assign QN = ~QP_aux;

endmodule